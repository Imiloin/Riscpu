module riscv (

    input wire clk,
    input wire rst,  // high is reset

    // inst_mem
    input  wire [31:0] inst_i,
    output wire [31:0] inst_addr_o,
    output wire        inst_ce_o,

    // data_mem
    input  wire [31:0] data_i,       // load data from data_mem
    output wire        data_we_o,
    output wire        data_ce_o,
    output wire [31:0] data_addr_o,
    output wire [31:0] data_o        // store data to data_mem

);

    // instance your module below





endmodule
