module IFID (
    input clk,
    input rst,
    input ifflush,  // flush the instruction, store a zero to IF/ID register