module MEM (  // Memory module, access the data memory
    input clk,
    input rst,
);

endmodule
